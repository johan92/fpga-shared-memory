import sm::*;

package sm_tb;

  `include "sm_cmd_driver.sv"
  `include "sm_res_monitor.sv"
  `include "sm_ref_model.sv"
  `include "sm_scoreboard.sv"

endpackage
